--
-- memif_def_sim.vhd - Simulation version of package 'memif_def'
--

package memif_def is

    constant memif_simulation : boolean := true;

end;

package body memif_def is

end;
