--
-- memif_def_synth.vhd - Synthesis version of package 'memif_def'
--

package memif_def is

    constant memif_simulation : boolean := false;

end;

package body memif_def is

end;
